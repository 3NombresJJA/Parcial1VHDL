  library IEEE;
use IEEE.std_logic_1164.all;

entity DivFreq is
	port
	(
		Clk	: in  std_logic;
		Sigue : in std_logic;
		out2 : buffer std_logic);
		
end DivFreq;

architecture Parque of DivFreq is

begin
ContadorSeg: process(clk)
variable count2 : integer range 0 to 25000000;
begin
	if(Sigue='1')then
		if (clk'event and clk='1') then
			count2 := count2 +1;
			if (count2 = 25000000) then 
				out2 <= not out2;
				count2 := 0;
			end if;
		end if;
	else
		out2<='0';
	end if;
end process;
end parque;