library verilog;
use verilog.vl_types.all;
entity ParcialV1_4_vlg_vec_tst is
end ParcialV1_4_vlg_vec_tst;
