library verilog;
use verilog.vl_types.all;
entity Cronometro_vlg_vec_tst is
end Cronometro_vlg_vec_tst;
