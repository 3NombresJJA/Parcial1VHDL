library verilog;
use verilog.vl_types.all;
entity ContadorenReversa_vlg_vec_tst is
end ContadorenReversa_vlg_vec_tst;
